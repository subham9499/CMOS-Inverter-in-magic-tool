* SPICE3 file created from inverter.ext - technology: scmos

.option scale=0.09u

M1000 out in vdd vdd pfet w=8 l=2
+  ad=40 pd=26 as=40 ps=26
M1001 out in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=20 ps=18
